netcdf domain_bci_fates_tutorial {
dimensions:
	nv = 4 ;
variables:
	double xc ;
		xc:_FillValue = NaN ;
		xc:long_name = "longitude of grid cell center" ;
		xc:units = "degrees_east" ;
		xc:bounds = "xv" ;
	double yc ;
		yc:_FillValue = NaN ;
		yc:long_name = "latitude of grid cell center" ;
		yc:units = "degrees_north" ;
		yc:bounds = "yv" ;
		yc:filter1 = " set_fv_pole_yc ON, yc = -+90 at j=1,j=nj" ;
	double xv(nv) ;
		xv:_FillValue = NaN ;
		xv:long_name = "longitude of grid cell verticies" ;
		xv:coordinates = "xc yc" ;
	double yv(nv) ;
		yv:_FillValue = NaN ;
		yv:long_name = "latitude of grid cell verticies" ;
		yv:coordinates = "xc yc" ;
	int mask ;
		mask:long_name = "domain mask" ;
		mask:note = "unitless" ;
		mask:comment = "0 value indicates cell is not active" ;
		mask:coordinates = "xc yc" ;
	double area ;
		area:_FillValue = NaN ;
		area:long_name = "area of grid cell in radians squared" ;
		area:units = "radian2" ;
		area:coordinates = "xc yc" ;
	double frac ;
		frac:_FillValue = NaN ;
		frac:coordinates = "xc yc" ;

// global attributes:
		:title = "CCSM domain data:" ;
		:Conventions = "CF-1.0" ;
		:source_code = "SVN $Id: gen_domain.F90 6671 2007-09-28 21:56:26Z kauff $" ;
		:SVN_url = " $URL: https://svn-ccsm-models.cgd.ucar.edu/tools/mapping/gen_domain/trunk/gen_domain.F90 $" ;
		:history = "created by kauff, 2009-02-06 12:19:29" ;
		:source = "/fis/cgd/cseg/csm/mapping/makemaps/fv1.9x2.5_gx1v6_090206/map_gx1v6_to_fv1.9x2.5_aave_da_090206.nc" ;
		:map_domain_a = "gx1v6, Present DP x1" ;
		:map_domain_b = "1.9x2.5 CAM finite volume grid" ;
		:map_grid_file_ocn = "/fis/cgd/cseg/csm/mapping/grids/gx1v6_090205.nc" ;
		:map_grid_file_atm = "/fis/cgd/cseg/csm/mapping/grids/fv1.9x2.5_060511.nc" ;
		:output_file1 = "domain.ocn.gx1v6.090206.nc" ;
		:output_file2 = "domain.lnd.fv1.9x2.5_gx1v6.090206.nc" ;
		:user_comment = "Standard CCSM3.1/4.0 domain specification file with fv pole fix" ;
data:

 xc = 280 ;

 yc = 8.5263157894736 ;

 xv = 278.75, 281.25, 281.25, 278.75 ;

 yv = 7.57894736842097, 7.57894736842097, 9.47368421052623, 9.47368421052623 ;

 mask = 1 ;

 area = 0.00142691220961584 ;

 frac = 1 ;
}
